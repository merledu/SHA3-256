`timescale 1ns / 1ps

module toptb();

        logic clk;
        logic rst;
        logic en;
       // logic [4:0] data_in; //5bit
       // logic [4:0] data_in; //8bit
        logic [39:0] data_in; //30bit
        //logic [1599:0] data_in; //1600bit
        logic [0:255] digest;
    
    Sha3_256 u_sha0 (
        .clk(clk),
        .rst(rst),
        .en(en),
        .datain(data_in),
        .digest(digest)
    );
    
    initial begin
    data_in = 40'h0;
//data_in = 40'h71696d6177;
//      data_in = 2320'h2E6E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D4148532E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;
        clk=1;
        rst=1;
        en=0;
        #2rst=0;
        #10data_in = 40'h1111111111;
        #10data_in = 40'h71696d6177;

        #2;
//        data_in = 2320'h2E6E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D4148532E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;

//        rst=0;
//        #10data_in = 40'h71696d6177;
//              data_in = 2320'h2E6E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D4148532E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;

        #20en=1;
        

      //  data_in=30'b1
; //5bit
     //  data_in = 1000'ha1b35c6e28f9d4723bc5817fa43d9e26b0e57fa2c68a14f77bcd3e6a58f10435be92d7b013f4a7c9256ebf8302917df85a1b03e5d489c2f67e18d4c76f3a59b24d2e9a7c134fb5789de4306a75b8c1023e5f9ab4c8d7e21bc75fa30147bd681efc97a524b8d6e35a21f7c0e93b5468c175da9e4b35cf037ab6e2d;
   
//   data_in = 40'h71696d6177;
//    data_in = 64'b0;
 //    DO    //  data_in = 1600'b1010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011;
 //   NOT    //  data_in = 1605'b000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011;
 //  CHANGE  //  data_in = 1630'b1000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011101000111010001110100011;
 // data_in = 4000'h2E737469622E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D4148532E737469622036353220332D616873206E6F20676E696B726F7720796C746E65727275632065726577206557202E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;
  // data_in = 2880'h2E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D4148532E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;
  // data_in = 1440'h2E796C696D616620332D4148532065687420666F2074726170207361202979676F6C6F6E6863655420646E612073647261646E61745320666F20657475746974736E49206C616E6F6974614E28205453494E2079622035313032206E692064657A69647261646E617473207361772074616874206E6F6974636E7566206873616820636968706172676F74707972632061207369202933206D687469726F676C412068736148206572756365532820332D414853;
    //data_in = 1600'b1110000010100101111001100001000101001010000110001111001100101111101100100111111111101111101010000001110000001000111110010111101000000110110110111011000010101011010001000010110010111010010111101001011110001010001010100001100110000100010111111010101001101000111100111000010010001111001111111011011110000111000110001110110100010000000000101100010010010011001011001100011010101110101101110111000101111001110011010110111000001010011111111011001100111100100101011001101100001110100101011101111111000111011100100000101000001011110001001011010100011001001100111110000101010011110110110111001101100110011101111100000100101010111111100100100110010010011011000111000010010110101100001110011100111000011101100000111000000100000000000100011101111010110110100001000101111001100111000110101010001110111100000110101001001010110011000100101111010100111001010111000011011101110000111010100001101011001111110000100101011101000010100000010010110000010101100101100110011011001011000010111101100101101110111110101111101111001110001000100111111110101001111110111100100000011011010111000111001001010000111000101011101001101111110001001111000110100111000101111101010100110111111100000101100010000111111100001011010100001100111111000111100111011000101111010010000010011001110000101101110001110010001010110000001011101010110001000010010000010010010000001100010111010000110000010001011101101010111011000011101100111101110100110111000011110001100011100000101001111110111011010001000100011100010100101101010110101010100111001010110101000000101000101100110011101111100111110010001101011110101110000111010011110010011011101011111101;
    //  data_in = 1600'hE0A5E6114A18F32FB27FEFA81C08F97A06DBB0AB442CBA5E978A2A19845FAA68F3848F3FB78718ED1002C4932CC6AEB77179CD6E0A7FB33C959B0E95DFC7720A0BC4B51933E153DB736677C12AFE49926C7096B0E738760E0400477ADA11799C6A8EF06A4ACC4BD4E570DDC3A86B3F095D0A04B056599B2C2F65BBEBEF3889FEA7EF206D71C9438AE9BF13C69C5F54DFC1621FC2D433F1E762F482670B71C8AC0BAB109049031743045DABB0ECF74DC3C63829FBB444714B56AA72B5028B33BE7C8D7AE1D3C9BAFD; 
  // data_in = 152'hfa71696D61777369656D616E796D6F6C6C6568;
 //  data_in = 5'b10011;
//data_in = 30'b011001011110110101100001010011;
   //data_in = 16'h9121;
      //  data_in = 1600'b1010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010;
       // data_in = 1600'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
      //  data_in = 16'habac;
     //data_in = 1600'ha3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3a3;
   //  data_in = 1600'hd8952d191b5363e97a476798995e23722e76de20d3629ace8a28e3cfefc51057999226ed23d6ae5c805f3fd0a8dfe19ff3d3763c15b7699034f6b2ec4d46af8ca864b980b3fc7697cfa81ff9e62352400e6bb69810a1973379cfdc6266c27288508854f1ef6609a8cb57937af747826f247d4107ffc043f0df35ea336b164a6246fac6c6b799f05467286757e733508062eccafb8360c6f9339e28f34f18767ac5ff6d593c9dfa8c2404ff227571373abd41c7518187971e25d2e8a53d9636348e2827ba4d2c6243;
     //  data_in = 1088'h24effea48fc3078fca8084c6881dbb9d944b0f3cc80797b4dda37631f5435cca47aa1101b2106f5f1bc8e3dbec9de63932a5f01f8c881a4a1c4733ffd61668902b7a7d5b8cbbbbbbbe5a2af29984846f004e95875aa8ff37e05bfcb375f27d5cff31df1d1a0616a634afa299e9172ac6ed46bd34adbaa05610386cf66308c001aca5b78e72b42562;
      //   data_in=2600'h2eba4b84dd377792ec6cd2e5a9a550684f2f112e28f91965043d82d90595780643c97878677f71564bb3ec72d0e0fbc7bba0a1649500be5987e26b8fcf028e5e5167d3f0c230c6c8d28c611822ef77e435a7e4b9f064588437aa6ec3b2253cce4cf581badfee9e2e78f4aedd151faa3c76e08c5d1ae5004d3a320c611bf6dc23be7e0863bc1358b709035f7e841ad751f33c3d6e4c283dae952c37b871f2c194e985e648f32f7313fdb29612b5309fea1c359f305544744b22158c565324effea48fc3078fca8084c6881dbb9d944b0f3cc80797b4dda37631f5435cca47aa1101b2106f5f1bc8e3dbec9de63932a5f01f8c881a4a1c4733ffd61668902b7a7d5b8cbbbbbbbe5a2af29984846f004e95875aa8ff37e05bfcb375f27d5cff31df1d1a0616a634afa299e9172ac6ed46bd34adbaa05610386cf66308c001aca5b78e72b42562; //8bit
     //  data_in=30'h197b5853; //30bit
         //data_in=1600'habcdefacdef; //1600bit
    
        #150;
        $finish;
    end
    
    always begin
            #2;
            clk = ~clk;
    end
    
    initial begin
            $dumpfile("sha.vcd");
            $dumpvars(0,toptb);
    end
    
endmodule
